// QsysCore.v

// Generated using ACDS version 13.0sp1 232 at 2020.06.09.07:20:42

`timescale 1 ps / 1 ps
module QsysCore (
		input  wire        clk_clk,                                                                                         //                                             clk.clk
		input  wire        reset_reset_n,                                                                                   //                                           reset.reset_n
		input  wire        spi_slave_to_avalon_mm_master_bridge_0_export_0_mosi_to_the_spislave_inst_for_spichain,          // spi_slave_to_avalon_mm_master_bridge_0_export_0.mosi_to_the_spislave_inst_for_spichain
		input  wire        spi_slave_to_avalon_mm_master_bridge_0_export_0_nss_to_the_spislave_inst_for_spichain,           //                                                .nss_to_the_spislave_inst_for_spichain
		inout  wire        spi_slave_to_avalon_mm_master_bridge_0_export_0_miso_to_and_from_the_spislave_inst_for_spichain, //                                                .miso_to_and_from_the_spislave_inst_for_spichain
		input  wire        spi_slave_to_avalon_mm_master_bridge_0_export_0_sclk_to_the_spislave_inst_for_spichain,          //                                                .sclk_to_the_spislave_inst_for_spichain
		output wire [31:0] pio_0_external_connection_export                                                                 //                       pio_0_external_connection.export
	);

	wire         spi_slave_to_avalon_mm_master_bridge_0_avalon_master_waitrequest;                                        // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:av_waitrequest -> spi_slave_to_avalon_mm_master_bridge_0:waitrequest_to_the_altera_avalon_packets_to_master_inst_for_spichain
	wire  [31:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_writedata;                                          // spi_slave_to_avalon_mm_master_bridge_0:writedata_from_the_altera_avalon_packets_to_master_inst_for_spichain -> spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:av_writedata
	wire  [31:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_address;                                            // spi_slave_to_avalon_mm_master_bridge_0:address_from_the_altera_avalon_packets_to_master_inst_for_spichain -> spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:av_address
	wire         spi_slave_to_avalon_mm_master_bridge_0_avalon_master_write;                                              // spi_slave_to_avalon_mm_master_bridge_0:write_from_the_altera_avalon_packets_to_master_inst_for_spichain -> spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:av_write
	wire         spi_slave_to_avalon_mm_master_bridge_0_avalon_master_read;                                               // spi_slave_to_avalon_mm_master_bridge_0:read_from_the_altera_avalon_packets_to_master_inst_for_spichain -> spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:av_read
	wire  [31:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdata;                                           // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:av_readdata -> spi_slave_to_avalon_mm_master_bridge_0:readdata_to_the_altera_avalon_packets_to_master_inst_for_spichain
	wire         spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdatavalid;                                      // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:av_readdatavalid -> spi_slave_to_avalon_mm_master_bridge_0:readdatavalid_to_the_altera_avalon_packets_to_master_inst_for_spichain
	wire   [3:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_byteenable;                                         // spi_slave_to_avalon_mm_master_bridge_0:byteenable_from_the_altera_avalon_packets_to_master_inst_for_spichain -> spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:av_byteenable
	wire         spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest;   // pio_0_s1_translator:uav_waitrequest -> spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_waitrequest
	wire   [2:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount;    // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_burstcount -> pio_0_s1_translator:uav_burstcount
	wire  [31:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_writedata;     // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_writedata -> pio_0_s1_translator:uav_writedata
	wire  [31:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_address;       // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_address -> pio_0_s1_translator:uav_address
	wire         spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_lock;          // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_lock -> pio_0_s1_translator:uav_lock
	wire         spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_write;         // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_write -> pio_0_s1_translator:uav_write
	wire         spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_read;          // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_read -> pio_0_s1_translator:uav_read
	wire  [31:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_readdata;      // pio_0_s1_translator:uav_readdata -> spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_readdata
	wire         spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess;   // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_debugaccess -> pio_0_s1_translator:uav_debugaccess
	wire   [3:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable;    // spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_byteenable -> pio_0_s1_translator:uav_byteenable
	wire         spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid; // pio_0_s1_translator:uav_readdatavalid -> spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:uav_readdatavalid
	wire  [31:0] pio_0_s1_translator_avalon_anti_slave_0_writedata;                                                       // pio_0_s1_translator:av_writedata -> pio_0:writedata
	wire   [1:0] pio_0_s1_translator_avalon_anti_slave_0_address;                                                         // pio_0_s1_translator:av_address -> pio_0:address
	wire         pio_0_s1_translator_avalon_anti_slave_0_chipselect;                                                      // pio_0_s1_translator:av_chipselect -> pio_0:chipselect
	wire         pio_0_s1_translator_avalon_anti_slave_0_write;                                                           // pio_0_s1_translator:av_write -> pio_0:write_n
	wire  [31:0] pio_0_s1_translator_avalon_anti_slave_0_readdata;                                                        // pio_0:readdata -> pio_0_s1_translator:av_readdata
	wire         rst_controller_reset_out_reset;                                                                          // rst_controller:reset_out -> [pio_0:reset_n, pio_0_s1_translator:reset, spi_slave_to_avalon_mm_master_bridge_0:reset_n, spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator:reset]

	SPISlaveToAvalonMasterBridge #(
		.SYNC_DEPTH (2)
	) spi_slave_to_avalon_mm_master_bridge_0 (
		.clk                                                                    (clk_clk),                                                                                         //           clk.clk
		.reset_n                                                                (~rst_controller_reset_out_reset),                                                                 //     clk_reset.reset_n
		.mosi_to_the_spislave_inst_for_spichain                                 (spi_slave_to_avalon_mm_master_bridge_0_export_0_mosi_to_the_spislave_inst_for_spichain),          //      export_0.export
		.nss_to_the_spislave_inst_for_spichain                                  (spi_slave_to_avalon_mm_master_bridge_0_export_0_nss_to_the_spislave_inst_for_spichain),           //              .export
		.miso_to_and_from_the_spislave_inst_for_spichain                        (spi_slave_to_avalon_mm_master_bridge_0_export_0_miso_to_and_from_the_spislave_inst_for_spichain), //              .export
		.sclk_to_the_spislave_inst_for_spichain                                 (spi_slave_to_avalon_mm_master_bridge_0_export_0_sclk_to_the_spislave_inst_for_spichain),          //              .export
		.address_from_the_altera_avalon_packets_to_master_inst_for_spichain     (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_address),                                    // avalon_master.address
		.byteenable_from_the_altera_avalon_packets_to_master_inst_for_spichain  (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_byteenable),                                 //              .byteenable
		.read_from_the_altera_avalon_packets_to_master_inst_for_spichain        (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_read),                                       //              .read
		.readdata_to_the_altera_avalon_packets_to_master_inst_for_spichain      (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdata),                                   //              .readdata
		.readdatavalid_to_the_altera_avalon_packets_to_master_inst_for_spichain (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdatavalid),                              //              .readdatavalid
		.waitrequest_to_the_altera_avalon_packets_to_master_inst_for_spichain   (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_waitrequest),                                //              .waitrequest
		.write_from_the_altera_avalon_packets_to_master_inst_for_spichain       (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_write),                                      //              .write
		.writedata_from_the_altera_avalon_packets_to_master_inst_for_spichain   (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_writedata)                                   //              .writedata
	);

	QsysCore_pio_0 pio_0 (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (pio_0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (pio_0_external_connection_export)                    // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator (
		.clk                      (clk_clk),                                                                                                 //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                          //                     reset.reset
		.uav_address              (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_byteenable),                                         //                          .byteenable
		.av_read                  (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_read),                                               //                          .read
		.av_readdata              (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_write),                                              //                          .write
		.av_writedata             (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                                                    //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                                    //               (terminated)
		.av_begintransfer         (1'b0),                                                                                                    //               (terminated)
		.av_chipselect            (1'b0),                                                                                                    //               (terminated)
		.av_lock                  (1'b0),                                                                                                    //               (terminated)
		.av_debugaccess           (1'b0),                                                                                                    //               (terminated)
		.uav_clken                (),                                                                                                        //               (terminated)
		.av_clken                 (1'b1),                                                                                                    //               (terminated)
		.uav_response             (2'b00),                                                                                                   //               (terminated)
		.av_response              (),                                                                                                        //               (terminated)
		.uav_writeresponserequest (),                                                                                                        //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                                    //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                                    //               (terminated)
		.av_writeresponsevalid    ()                                                                                                         //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_0_s1_translator (
		.clk                      (clk_clk),                                                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                          //                    reset.reset
		.uav_address              (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read                 (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write                (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest          (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata             (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata            (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock                 (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess          (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address               (pio_0_s1_translator_avalon_anti_slave_0_address),                                                         //      avalon_anti_slave_0.address
		.av_write                 (pio_0_s1_translator_avalon_anti_slave_0_write),                                                           //                         .write
		.av_readdata              (pio_0_s1_translator_avalon_anti_slave_0_readdata),                                                        //                         .readdata
		.av_writedata             (pio_0_s1_translator_avalon_anti_slave_0_writedata),                                                       //                         .writedata
		.av_chipselect            (pio_0_s1_translator_avalon_anti_slave_0_chipselect),                                                      //                         .chipselect
		.av_read                  (),                                                                                                        //              (terminated)
		.av_begintransfer         (),                                                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                                                        //              (terminated)
		.av_burstcount            (),                                                                                                        //              (terminated)
		.av_byteenable            (),                                                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                                        //              (terminated)
		.av_lock                  (),                                                                                                        //              (terminated)
		.av_clken                 (),                                                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                                                    //              (terminated)
		.av_debugaccess           (),                                                                                                        //              (terminated)
		.av_outputenable          (),                                                                                                        //              (terminated)
		.uav_response             (),                                                                                                        //              (terminated)
		.av_response              (2'b00),                                                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                     //              (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
